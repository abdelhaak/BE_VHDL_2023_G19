
module avaloon_cmps (
	avalon_cpt_0_conduit_end_beginbursttransfer,
	clk_clk);	

	input		avalon_cpt_0_conduit_end_beginbursttransfer;
	input		clk_clk;
endmodule
