library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity avaloon_verin is
port ( 	clk, chipselect, write_n, reset_n: in std_logic;
			writedata : in std_logic_vector (31 downto 0);
			address: std_logic_vector (3 downto 0);
			readdata : out std_logic_vector (31 downto 0);
			out_pwm : out std_logic;
			out_sens : out std_logic;
			cs : out std_logic
			);
end avaloon_verin;

architecture bhv of avaloon_verin is
---- Declaration des signaux

  signal s_freq, s_duty, s_bg, s_bd : std_logic_vector (15 downto 0);
  signal s_config : std_logic_vector (4 downto 0);
  signal raz_n, enable_pwm, sens :  std_logic;
  signal angle_barre :  std_logic_vector (11 downto 0);
  signal butee_d, butee_g, freq, duty : std_logic_vector (15 downto 0);
  signal fd, fg: std_logic;
  signal clk_1M, clk_50, data_in, enable, f_g, f_d : std_logic;
  signal data_out: std_logic_vector (11 downto 0);




----- COMPOSANT gestion_pwm
COMPONENT gestion_pwm
	PORT(
	clk_50Mhz, reset_n : in std_logic;
	freq, duty : in std_logic_vector (15 downto 0);
	out_pwm_sig : out std_logic
		 );
END COMPONENT;


----- COMPOSANT fct_mcp3201

COMPONENT fct_mcp
	PORT(
	clk_50Mhz : in std_logic;
	raz_n : in std_logic;
	data_in : in std_logic;
	clk_adc : out std_logic;
	cs_out : out std_logic;
	data_out : out std_logic_vector(11 downto 0)
		 );
END COMPONENT;



----- COMPOSANT control_butee
COMPONENT control_butee
	PORT(
	pwm_in, sens, enable: in std_logic;
	butee_g, butee_d : in std_logic_vector (15 downto 0);
	angle_barre : in std_logic_vector (11 downto 0);
	out_pwm, out_sens, f_g, f_d : out std_logic
		 );
END COMPONENT;

signal pwm_wire : std_logic;
signal angle_barre_wire :std_logic_vector(11 downto 0);

begin 
data_out <= angle_barre_wire;




------ POrt map de gestion pwm
bbv_inst1 : gestion_pwm 
port map(
		 clk_50Mhz => clk_50,
		 reset_n => reset_n,
		 duty => duty,
		 freq => freq,
		 out_pwm_sig => pwm_wire
			);



------ POrt map de fct_mcp	
bbv_inst2 : fct_mcp
port map(
			clk_50Mhz  => clk_50,
			raz_n   => raz_n, 
			data_in => data_in, 
			clk_adc  => clk_1M, 
			cs_out   => cs, 
			data_out=> angle_barre_wire
			);
			

------ POrt map de control_butee	

bbv_inst3 : control_butee 
port map(
	    pwm_in => pwm_wire,
		 sens => sens,
		 enable => enable,
		 angle_barre => angle_barre_wire,
		 butee_d => butee_d,
		 butee_g => butee_g,
		 out_pwm => out_pwm,
		 out_sens => out_sens,
		 f_g => f_g ,
		 f_d => f_d
		 );
		
	
	
process_write: process (clk, reset_n)
begin
	if reset_n = '0' then
		freq <= (others => '0');
		duty <= (others => '0');
		s_config <= (others => '0');
		butee_g <= (others => '0');
		butee_d <= (others => '0');
	elsif clk'event and clk = '1' then
		if chipselect ='1' and write_n = '0' then
			if address = "0000" then
				freq <= writedata(15 downto 0);
				s_freq <=  writedata(15 downto 0);
				duty <= writedata(31 downto 16);
				s_duty <=  writedata(31 downto 16);
			end if;
			if address = "0001" then
				butee_g <= writedata (15 downto 0);
				s_bg <=  writedata(15 downto 0);
				butee_d <= writedata (31 downto 16);
				s_bd <=  writedata(31 downto 16);
			end if;
			if address = "0010" then
				s_config(2 downto 0) <=  writedata(2 downto 0);
				s_config(3) <= fd;
				s_config(4) <= fg;
				raz_n <= s_config(0);
				enable_pwm <= s_config(1);
				sens <= s_config(2);

		end if;
	end if;
  end if;
end process process_write;
  
  
process_Read:process (address, angle_barre, s_freq, s_duty, s_bg, s_bd, s_config)

begin

	case address is
		when "0000" => readdata <= s_duty & s_freq ;
		when "0001" => readdata <= s_bd & s_bg ;
		when "0010" => readdata <= "000000000000000000000000000" & s_config ;
		when "0101" => readdata <= "00000000000000000000" & angle_barre ;
		when others => readdata <= (others => '0');
	end case;

END PROCESS process_Read ;
	
end bhv;