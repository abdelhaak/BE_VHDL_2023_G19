
module avalon_cpt (
	clk_clk,
	cs_writeresponsevalid_n,
	out_pwm_writeresponsevalid_n,
	out_sens_writeresponsevalid_n);	

	input		clk_clk;
	output		cs_writeresponsevalid_n;
	output		out_pwm_writeresponsevalid_n;
	output		out_sens_writeresponsevalid_n;
endmodule
